
module RoundFunction(a,
                     key0,
                     key2,
                     rc,
                     sbox_type,
                     b);

input [127:0] a;
input [31:0] key0;
input [31:0] key2;
input [5:0]  rc;
input        sbox_type;
output[127:0] b;

// ------------------------------

wire [31:0] a0,a1,a2,a3;
wire [31:0] s0,s1,s2,s3;
wire [31:0] p0,p1,p2,p3;
wire [31:0] b0,b1,b2,b3;

// ------------------------------

assign a0 = {a[124],a[120],a[116],a[112],a[108],a[104],a[100],a[96],a[92],a[88],a[84],a[80],a[76],a[72],a[68],a[64],a[60],a[56],a[52],a[48],a[44],a[40],a[36],a[32],a[28],a[24],a[20],a[16],a[12],a[8],a[4],a[0] };
assign a1 = {a[125],a[121],a[117],a[113],a[109],a[105],a[101],a[97],a[93],a[89],a[85],a[81],a[77],a[73],a[69],a[65],a[61],a[57],a[53],a[49],a[45],a[41],a[37],a[33],a[29],a[25],a[21],a[17],a[13],a[9],a[5],a[1] };
assign a2 = {a[126],a[122],a[118],a[114],a[110],a[106],a[102],a[98],a[94],a[90],a[86],a[82],a[78],a[74],a[70],a[66],a[62],a[58],a[54],a[50],a[46],a[42],a[38],a[34],a[30],a[26],a[22],a[18],a[14],a[10],a[6],a[2]};
assign a3 = {a[127],a[123],a[119],a[115],a[111],a[107],a[103],a[99],a[95],a[91],a[87],a[83],a[79],a[75],a[71],a[67],a[63],a[59],a[55],a[51],a[47],a[43],a[39],a[35],a[31],a[27],a[23],a[19],a[15],a[11],a[7],a[3]};

// ------------------------------
SubCells sc0(a0,a1,a2,a3,
             sbox_type,
             s0,s1,s2,s3);

PermBits pm0(s0,s1,s2,s3,
             p0,p1,p2,p3);

AddRoundKey ak0(p0,p1,p2,p3,
                key0,
                key2,
                rc,
                b0,b1,b2,b3);

// ------------------------------

assign b={b3[31],b2[31],b1[31],b0[31],
          b3[30],b2[30],b1[30],b0[30],
          b3[29],b2[29],b1[29],b0[29], 
          b3[28],b2[28],b1[28],b0[28], 
          b3[27],b2[27],b1[27],b0[27], 
          b3[26],b2[26],b1[26],b0[26], 
          b3[25],b2[25],b1[25],b0[25],
          b3[24],b2[24],b1[24],b0[24],
          b3[23],b2[23],b1[23],b0[23],
          b3[22],b2[22],b1[22],b0[22],
          b3[21],b2[21],b1[21],b0[21],
          b3[20],b2[20],b1[20],b0[20],
          b3[19],b2[19],b1[19],b0[19], 
          b3[18],b2[18],b1[18],b0[18], 
          b3[17],b2[17],b1[17],b0[17], 
          b3[16],b2[16],b1[16],b0[16], 
          b3[15],b2[15],b1[15],b0[15],
          b3[14],b2[14],b1[14],b0[14],
          b3[13],b2[13],b1[13],b0[13],
          b3[12],b2[12],b1[12],b0[12],
          b3[11],b2[11],b1[11],b0[11],
          b3[10],b2[10],b1[10],b0[10],
          b3[9] ,b2[9] ,b1[9] ,b0[9] ,
          b3[8] ,b2[8] ,b1[8] ,b0[8] ,
          b3[7] ,b2[7] ,b1[7] ,b0[7] ,
          b3[6] ,b2[6] ,b1[6] ,b0[6] ,
          b3[5] ,b2[5] ,b1[5] ,b0[5] ,
          b3[4] ,b2[4] ,b1[4] ,b0[4] ,
          b3[3] ,b2[3] ,b1[3] ,b0[3] ,
          b3[2] ,b2[2] ,b1[2] ,b0[2] ,
          b3[1] ,b2[1] ,b1[1] ,b0[1] ,
          b3[0] ,b2[0] ,b1[0] ,b0[0] };

endmodule


