
module RoundFunction(a,
                     key,
                     rc,
                     sbox_type,
                     b);

input [63:0] a;
input [31:0] key;
input [5:0]  rc;
input        sbox_type;
output[63:0] b;

// ------------------------------

wire [15:0] a0,a1,a2,a3;
wire [15:0] s0,s1,s2,s3;
wire [15:0] p0,p1,p2,p3;
wire [15:0] b0,b1,b2,b3;

// ------------------------------

assign a0 = {a[60],a[56],a[52],a[48],a[44],a[40],a[36],a[32],a[28],a[24],a[20],a[16],a[12],a[8] ,a[4],a[0]};
assign a1 = {a[61],a[57],a[53],a[49],a[45],a[41],a[37],a[33],a[29],a[25],a[21],a[17],a[13],a[9] ,a[5],a[1]};
assign a2 = {a[62],a[58],a[54],a[50],a[46],a[42],a[38],a[34],a[30],a[26],a[22],a[18],a[14],a[10],a[6],a[2]};
assign a3 = {a[63],a[59],a[55],a[51],a[47],a[43],a[39],a[35],a[31],a[27],a[23],a[19],a[15],a[11],a[7],a[3]};

// ------------------------------
SubCells sc0(a0,a1,a2,a3,
             sbox_type,
             s0,s1,s2,s3);

PermBits pm0(s0,s1,s2,s3,
             p0,p1,p2,p3);

AddRoundKey ak0(p0,p1,p2,p3,
                key,
                rc,
                b0,b1,b2,b3);

// ------------------------------

assign b={b3[15],b2[15],b1[15],b0[15],
          b3[14],b2[14],b1[14],b0[14],
          b3[13],b2[13],b1[13],b0[13],
          b3[12],b2[12],b1[12],b0[12],
          b3[11],b2[11],b1[11],b0[11],
          b3[10],b2[10],b1[10],b0[10],
          b3[9] ,b2[9] ,b1[9] ,b0[9] ,
          b3[8] ,b2[8] ,b1[8] ,b0[8] ,
          b3[7] ,b2[7] ,b1[7] ,b0[7] ,
          b3[6] ,b2[6] ,b1[6] ,b0[6] ,
          b3[5] ,b2[5] ,b1[5] ,b0[5] ,
          b3[4] ,b2[4] ,b1[4] ,b0[4] ,
          b3[3] ,b2[3] ,b1[3] ,b0[3] ,
          b3[2] ,b2[2] ,b1[2] ,b0[2] ,
          b3[1] ,b2[1] ,b1[1] ,b0[1] ,
          b3[0] ,b2[0] ,b1[0] ,b0[0] };

endmodule