
module PermBits(a0,a1,a2,a3,
                b0,b1,b2,b3);

input [31:0] a0,a1,a2,a3;
output[31:0] b0,b1,b2,b3;

assign b0[0] = a0[0];
assign b0[24] = a0[1];
assign b0[16] = a0[2];
assign b0[8] = a0[3];
assign b0[1] = a0[4];
assign b0[25] = a0[5];
assign b0[17] = a0[6];
assign b0[9] = a0[7];
assign b0[2] = a0[8];
assign b0[26] = a0[9];
assign b0[18] = a0[10];
assign b0[10] = a0[11];
assign b0[3] = a0[12];
assign b0[27] = a0[13];
assign b0[19] = a0[14];
assign b0[11] = a0[15];
assign b0[4] = a0[16];
assign b0[28] = a0[17];
assign b0[20] = a0[18];
assign b0[12] = a0[19];
assign b0[5] = a0[20];
assign b0[29] = a0[21];
assign b0[21] = a0[22];
assign b0[13] = a0[23];
assign b0[6] = a0[24];
assign b0[30] = a0[25];
assign b0[22] = a0[26];
assign b0[14] = a0[27];
assign b0[7] = a0[28];
assign b0[31] = a0[29];
assign b0[23] = a0[30];
assign b0[15] = a0[31];
assign b1[8] = a1[0];
assign b1[0] = a1[1];
assign b1[24] = a1[2];
assign b1[16] = a1[3];
assign b1[9] = a1[4];
assign b1[1] = a1[5];
assign b1[25] = a1[6];
assign b1[17] = a1[7];
assign b1[10] = a1[8];
assign b1[2] = a1[9];
assign b1[26] = a1[10];
assign b1[18] = a1[11];
assign b1[11] = a1[12];
assign b1[3] = a1[13];
assign b1[27] = a1[14];
assign b1[19] = a1[15];
assign b1[12] = a1[16];
assign b1[4] = a1[17];
assign b1[28] = a1[18];
assign b1[20] = a1[19];
assign b1[13] = a1[20];
assign b1[5] = a1[21];
assign b1[29] = a1[22];
assign b1[21] = a1[23];
assign b1[14] = a1[24];
assign b1[6] = a1[25];
assign b1[30] = a1[26];
assign b1[22] = a1[27];
assign b1[15] = a1[28];
assign b1[7] = a1[29];
assign b1[31] = a1[30];
assign b1[23] = a1[31];
assign b2[16] = a2[0];
assign b2[8] = a2[1];
assign b2[0] = a2[2];
assign b2[24] = a2[3];
assign b2[17] = a2[4];
assign b2[9] = a2[5];
assign b2[1] = a2[6];
assign b2[25] = a2[7];
assign b2[18] = a2[8];
assign b2[10] = a2[9];
assign b2[2] = a2[10];
assign b2[26] = a2[11];
assign b2[19] = a2[12];
assign b2[11] = a2[13];
assign b2[3] = a2[14];
assign b2[27] = a2[15];
assign b2[20] = a2[16];
assign b2[12] = a2[17];
assign b2[4] = a2[18];
assign b2[28] = a2[19];
assign b2[21] = a2[20];
assign b2[13] = a2[21];
assign b2[5] = a2[22];
assign b2[29] = a2[23];
assign b2[22] = a2[24];
assign b2[14] = a2[25];
assign b2[6] = a2[26];
assign b2[30] = a2[27];
assign b2[23] = a2[28];
assign b2[15] = a2[29];
assign b2[7] = a2[30];
assign b2[31] = a2[31];
assign b3[24] = a3[0];
assign b3[16] = a3[1];
assign b3[8] = a3[2];
assign b3[0] = a3[3];
assign b3[25] = a3[4];
assign b3[17] = a3[5];
assign b3[9] = a3[6];
assign b3[1] = a3[7];
assign b3[26] = a3[8];
assign b3[18] = a3[9];
assign b3[10] = a3[10];
assign b3[2] = a3[11];
assign b3[27] = a3[12];
assign b3[19] = a3[13];
assign b3[11] = a3[14];
assign b3[3] = a3[15];
assign b3[28] = a3[16];
assign b3[20] = a3[17];
assign b3[12] = a3[18];
assign b3[4] = a3[19];
assign b3[29] = a3[20];
assign b3[21] = a3[21];
assign b3[13] = a3[22];
assign b3[5] = a3[23];
assign b3[30] = a3[24];
assign b3[22] = a3[25];
assign b3[14] = a3[26];
assign b3[6] = a3[27];
assign b3[31] = a3[28];
assign b3[23] = a3[29];
assign b3[15] = a3[30];
assign b3[7] = a3[31];

endmodule